module sensorpro

fn main() {
}
